module ControlUnit (
);
endmodule