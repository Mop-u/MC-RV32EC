module TagMgmt_Testbench ();
initial $finish();

endmodule